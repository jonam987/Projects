typedef uvm_sequencer#(rd_tx) read_sqr;
